`include "dpu.v"

module shape (clk, rst, xin, yin, xout, yout);
   input clk, rst;
   wire clk, rst;
   input signed [31:0] xin;
   input signed [31:0] yin;
   output signed [31:0] xout;
   output signed [31:0] yout;

   wire signed [31:0]   xin;
   wire signed [31:0]   yin;

   wire signed [31:0]   xout;
   wire signed [31:0]   yout;

   wire signed [31:0]   xout1;
   wire signed [31:0]   xout2;
   wire signed [31:0]   xout3;
   wire signed [31:0]   xout4;
   wire signed [31:0]   xout5;
   wire signed [31:0]   xout6;
   wire signed [31:0]   xout7;
   wire signed [31:0]   xout8;
   wire signed [31:0]   xout9;
   wire signed [31:0]   xout10;
   wire signed [31:0]   xout11;
   wire signed [31:0]   xout12;
   wire signed [31:0]   xout13;
   wire signed [31:0]   xout14;
   wire signed [31:0]   xout15;
   wire signed [31:0]   xout16;
   wire signed [31:0]   xout17;
   wire signed [31:0]   xout18;
   wire signed [31:0]   xout19;
   wire signed [31:0]   xout20;
   wire signed [31:0]   xout21;
   wire signed [31:0]   xout22;
   wire signed [31:0]   xout23;
   wire signed [31:0]   xout24;
   wire signed [31:0]   xout25;
   wire signed [31:0]   xout26;
   wire signed [31:0]   xout27;
   wire signed [31:0]   xout28;
   wire signed [31:0]   xout29;
   wire signed [31:0]   xout30;
   wire signed [31:0]   xout31;
   wire signed [31:0]   xout32;

   wire signed [31:0]   yout1;
   wire signed [31:0]   yout2;
   wire signed [31:0]   yout3;
   wire signed [31:0]   yout4;
   wire signed [31:0]   yout5;
   wire signed [31:0]   yout6;
   wire signed [31:0]   yout7;
   wire signed [31:0]   yout8;
   wire signed [31:0]   yout9;
   wire signed [31:0]   yout10;
   wire signed [31:0]   yout11;
   wire signed [31:0]   yout12;
   wire signed [31:0]   yout13;
   wire signed [31:0]   yout14;
   wire signed [31:0]   yout15;
   wire signed [31:0]   yout16;
   wire signed [31:0]   yout17;
   wire signed [31:0]   yout18;
   wire signed [31:0]   yout19;
   wire signed [31:0]   yout20;
   wire signed [31:0]   yout21;
   wire signed [31:0]   yout22;
   wire signed [31:0]   yout23;
   wire signed [31:0]   yout24;
   wire signed [31:0]   yout25;
   wire signed [31:0]   yout26;
   wire signed [31:0]   yout27;
   wire signed [31:0]   yout28;
   wire signed [31:0]   yout29;
   wire signed [31:0]   yout30;
   wire signed [31:0]   yout31;
   wire signed [31:0]   yout32;

   localparam w1 = 32'sd1235;
   localparam w2 = 32'sd115;
   localparam w3 = -32'sd1280;
   localparam w4 = -32'sd2732;
   localparam w5 = -32'sd3965;
   localparam w6 = -32'sd4686;
   localparam w7 = -32'sd4627;
   localparam w8 = -32'sd3592;
   localparam w9 = -32'sd1496;
   localparam w10 = 32'sd1612;
   localparam w11 = 32'sd5538;
   localparam w12 = 32'sd9964;
   localparam w13 = 32'sd14478;
   localparam w14 = 32'sd18623;
   localparam w15 = 32'sd21960;
   localparam w16 = 32'sd24125;
   localparam w17 = 32'sd24874;
   localparam w18 = 32'sd24125;
   localparam w19 = 32'sd21960;
   localparam w20 = 32'sd18623;
   localparam w21 = 32'sd14478;
   localparam w22 = 32'sd9964;
   localparam w23 = 32'sd5538;
   localparam w24 = 32'sd1612;
   localparam w25 = -32'sd1496;
   localparam w26 = -32'sd3592;
   localparam w27 = -32'sd4627;
   localparam w28 = -32'sd4686;
   localparam w29 = -32'sd3965;
   localparam w30 = -32'sd2732;
   localparam w31 = -32'sd1280;
   localparam w32 = 32'sd115;
   localparam w33 = 32'sd1235;

   dpu stage1 ( .clk(clk), .rst(rst), .w(w1), .xin(xin), .yin(yin), .xout(xout1), .yout(yout1) );
   dpu stage2 ( .clk(clk), .rst(rst), .w(w2), .xin(xout1), .yin(yout1), .xout(xout2), .yout(yout2) );
   dpu stage3 ( .clk(clk), .rst(rst), .w(w3), .xin(xout2), .yin(yout2), .xout(xout3), .yout(yout3) );
   dpu stage4 ( .clk(clk), .rst(rst), .w(w4), .xin(xout3), .yin(yout3), .xout(xout4), .yout(yout4) );
   dpu stage5 ( .clk(clk), .rst(rst), .w(w5), .xin(xout4), .yin(yout4), .xout(xout5), .yout(yout5) );
   dpu stage6 ( .clk(clk), .rst(rst), .w(w6), .xin(xout5), .yin(yout5), .xout(xout6), .yout(yout6) );
   dpu stage7 ( .clk(clk), .rst(rst), .w(w7), .xin(xout6), .yin(yout6), .xout(xout7), .yout(yout7) );
   dpu stage8 ( .clk(clk), .rst(rst), .w(w8), .xin(xout7), .yin(yout7), .xout(xout8), .yout(yout8) );
   dpu stage9 ( .clk(clk), .rst(rst), .w(w9), .xin(xout8), .yin(yout8), .xout(xout9), .yout(yout9) );
   dpu stage10 ( .clk(clk), .rst(rst), .w(w10), .xin(xout9), .yin(yout9), .xout(xout10), .yout(yout10) );
   dpu stage11 ( .clk(clk), .rst(rst), .w(w11), .xin(xout10), .yin(yout10), .xout(xout11), .yout(yout11) );
   dpu stage12 ( .clk(clk), .rst(rst), .w(w12), .xin(xout11), .yin(yout11), .xout(xout12), .yout(yout12) );
   dpu stage13 ( .clk(clk), .rst(rst), .w(w13), .xin(xout12), .yin(yout12), .xout(xout13), .yout(yout13) );
   dpu stage14 ( .clk(clk), .rst(rst), .w(w14), .xin(xout13), .yin(yout13), .xout(xout14), .yout(yout14) );
   dpu stage15 ( .clk(clk), .rst(rst), .w(w15), .xin(xout14), .yin(yout14), .xout(xout15), .yout(yout15) );
   dpu stage16 ( .clk(clk), .rst(rst), .w(w16), .xin(xout15), .yin(yout15), .xout(xout16), .yout(yout16) );
   dpu stage17 ( .clk(clk), .rst(rst), .w(w17), .xin(xout16), .yin(yout16), .xout(xout17), .yout(yout17) );
   dpu stage18 ( .clk(clk), .rst(rst), .w(w18), .xin(xout17), .yin(yout17), .xout(xout18), .yout(yout18) );
   dpu stage19 ( .clk(clk), .rst(rst), .w(w19), .xin(xout18), .yin(yout18), .xout(xout19), .yout(yout19) );
   dpu stage20 ( .clk(clk), .rst(rst), .w(w20), .xin(xout19), .yin(yout19), .xout(xout20), .yout(yout20) );
   dpu stage21 ( .clk(clk), .rst(rst), .w(w21), .xin(xout20), .yin(yout20), .xout(xout21), .yout(yout21) );
   dpu stage22 ( .clk(clk), .rst(rst), .w(w22), .xin(xout21), .yin(yout21), .xout(xout22), .yout(yout22) );
   dpu stage23 ( .clk(clk), .rst(rst), .w(w23), .xin(xout22), .yin(yout22), .xout(xout23), .yout(yout23) );
   dpu stage24 ( .clk(clk), .rst(rst), .w(w24), .xin(xout23), .yin(yout23), .xout(xout24), .yout(yout24) );
   dpu stage25 ( .clk(clk), .rst(rst), .w(w25), .xin(xout24), .yin(yout24), .xout(xout25), .yout(yout25) );
   dpu stage26 ( .clk(clk), .rst(rst), .w(w26), .xin(xout25), .yin(yout25), .xout(xout26), .yout(yout26) );
   dpu stage27 ( .clk(clk), .rst(rst), .w(w27), .xin(xout26), .yin(yout26), .xout(xout27), .yout(yout27) );
   dpu stage28 ( .clk(clk), .rst(rst), .w(w28), .xin(xout27), .yin(yout27), .xout(xout28), .yout(yout28) );
   dpu stage29 ( .clk(clk), .rst(rst), .w(w29), .xin(xout28), .yin(yout28), .xout(xout29), .yout(yout29) );
   dpu stage30 ( .clk(clk), .rst(rst), .w(w30), .xin(xout29), .yin(yout29), .xout(xout30), .yout(yout30) );
   dpu stage31 ( .clk(clk), .rst(rst), .w(w31), .xin(xout30), .yin(yout30), .xout(xout31), .yout(yout31) );
   dpu stage32 ( .clk(clk), .rst(rst), .w(w32), .xin(xout31), .yin(yout31), .xout(xout32), .yout(yout32) );
   dpu stage33 ( .clk(clk), .rst(rst), .w(w33), .xin(xout32), .yin(yout32), .xout(xout), .yout(yout) );
endmodule
